grammar edu:umn:cs:melt:exts:ableC:exponent;

exports edu:umn:cs:melt:exts:ableC:exponent:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:exponent:concretesyntax;